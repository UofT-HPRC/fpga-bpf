//Copyright 2020 Marco Merlini. This file is part of the fpga-bpf project,
//whose license information can be found at 
//https://github.com/UofT-HPRC/fpga-bpf/blob/master/LICENSE

`timescale 1ns / 1ps

/*

module_template.v

Replace innards with desired logic

*/

module module_template # (
    parameter X = 5
) (
    input wire clk,
    input wire rst
    
    //...
);
    /************************************/
    /**Forward-declare internal signals**/
    /************************************/
    
    
    
    /***************************************/
    /**Assign internal signals from inputs**/
    /***************************************/
    
    
    
    /************************************/
    /**Helpful names for neatening code**/
    /************************************/
    
    
    
    /****************/
    /**Do the logic**/
    /****************/
    
    
    
    /****************************************/
    /**Assign outputs from internal signals**/
    /****************************************/



endmodule
