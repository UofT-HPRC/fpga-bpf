`timescale 1ns / 1ps

/*

module_template.v

Replace innards with desired logic

*/

module module_template # (
    parameter X = Y
) (
    input wire clk,
    input wire rst,
    
    ...
);

    //Code here

endmodule
