`timescale 1ns / 1ps

`include "p3.v"

module p3_tb;




endmodule
