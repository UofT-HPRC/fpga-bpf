`timescale 1ns / 1ps

/*

module_template.v

Replace innards with desired logic

*/

module module_template # (
    parameter X = Y
) (
    input wire clk,
    input wire rst,
    
    ...
);
    /************************************/
    /**Forward-declare internal signals**/
    /************************************/
    
    
    
    /***************************************/
    /**Assign internal signals from inputs**/
    /***************************************/
    
    
    
    /************************************/
    /**Helpful names for neatening code**/
    /************************************/
    
    
    
    /****************/
    /**Do the logic**/
    /****************/
    
    
    
    /****************************************/
    /**Assign outputs from internal signals**/
    /****************************************/



endmodule
